entity tb is
end tb;

architecture bench of tb is

	--COMPONENTES
	

	--SINAIS
	

	--for DESL_LEFT : SHFTL use entity work.SHFTL;

	begin

	--DESL_LEFT : SHFTL port map (I => A, S => SEL, Y => F);


	process
	begin
		


		wait;
		end process;

end bench;

