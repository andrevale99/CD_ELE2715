--==============================================================================================
--				LOGICA DO SUBTRATOR COMPLETO
--==============================================================================================