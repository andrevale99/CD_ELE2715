entity ckt_tb is
end ckt_tb;
	
architecture bench of ckt_tb is
	
	begin
		
	
	process
	begin
		
		wait;
	end process;

end bench;