--===========================================================
-- MUX ARRAY 10 BITS INPUT COM 3 BITS DE SELECAO
--===========================================================

entity MUX13B4S is
	port ( I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16 : in bit_vector(12 downto 0);
			S : in bit_vector(3 downto 0);
			Q : out bit_vector(12 downto 0));
end MUX13B4S;

architecture ckt of MUX13B4S is

    component MUX4S is
        port ( I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16 : in bit;
                S : in bit_vector(3 downto 0);
                Q : out bit);
    end component;

begin 

		Q1 : MUX4S port map ( I1(0), I2(0),  I3(0),  I4(0),  I5(0),  I6(0),  I7(0),  I8(0),  I9(0),  I10(0),  I11(0),  I12(0),  I13(0),  I14(0),  I15(0),  I16(0),  S, Q(0));
		Q2 : MUX4S port map ( I1(1), I2(1),  I3(1),  I4(1),  I5(1),  I6(1),  I7(1),  I8(1),  I9(1),  I10(1),  I11(1),  I12(1),  I13(1),  I14(1),  I15(1),  I16(1),  S, Q(1));
		Q3 : MUX4S port map ( I1(2), I2(2),  I3(2),  I4(2),  I5(2),  I6(2),  I7(2),  I8(2),  I9(2),  I10(2),  I11(2),  I12(2),  I13(2),  I14(2),  I15(2),  I16(2),  S, Q(2));
		Q4 : MUX4S port map ( I1(3), I2(3),  I3(3),  I4(3),  I5(3),  I6(3),  I7(3),  I8(3),  I9(3),  I10(3),  I11(3),  I12(3),  I13(3),  I14(3),  I15(3),  I16(3),  S, Q(3));
		Q5 : MUX4S port map ( I1(4), I2(4),  I3(4),  I4(4),  I5(4),  I6(4),  I7(4),  I8(4),  I9(4),  I10(4),  I11(4),  I12(4),  I13(4),  I14(4),  I15(4),  I16(4),  S, Q(4));
		Q6 : MUX4S port map ( I1(5), I2(5),  I3(5),  I4(5),  I5(5),  I6(5),  I7(5),  I8(5),  I9(5),  I10(5),  I11(5),  I12(5),  I13(5),  I14(5),  I15(5),  I16(5),  S, Q(5));
		Q7 : MUX4S port map ( I1(6), I2(6),  I3(6),  I4(6),  I5(6),  I6(6),  I7(6),  I8(6),  I9(6),  I10(6),  I11(6),  I12(6),  I13(6),  I14(6),  I15(6),  I16(6),  S, Q(6));
		Q8 : MUX4S port map ( I1(7), I2(7),  I3(7),  I4(7),  I5(7),  I6(7),  I7(7),  I8(7),  I9(7),  I10(7),  I11(7),  I12(7),  I13(7),  I14(7),  I15(7),  I16(7),  S, Q(7));
		Q9 : MUX4S port map ( I1(8), I2(8),  I3(8),  I4(8),  I5(8),  I6(8),  I7(8),  I8(8),  I9(8),  I10(8),  I11(8),  I12(8),  I13(8),  I14(8),  I15(8),  I16(8),  S, Q(8));
	   Q10 : MUX4S port map ( I1(9), I2(9),  I3(9),  I4(9),  I5(9),  I6(9),  I7(9),  I8(9),  I9(9),  I10(9),  I11(9),  I12(9),  I13(9),  I14(9),  I15(9),  I16(9),  S, Q(9));
       Q11 : MUX4S port map (I1(10), I2(10), I3(10), I4(10), I5(10), I6(10), I7(10), I8(10), I9(10), I10(10), I11(10), I12(10), I13(10), I14(10), I15(10), I16(10), S, Q(10));
       Q12 : MUX4S port map (I1(11), I2(11), I3(11), I4(11), I5(11), I6(11), I7(11), I8(11), I9(11), I10(11), I11(11), I12(11), I13(11), I14(11), I15(11), I16(11), S, Q(11));
       Q13 : MUX4S port map (I1(12), I2(12), I3(12), I4(12), I5(12), I6(12), I7(12), I8(12), I9(12), I10(12), I11(12), I12(12), I13(12), I14(12), I15(12), I16(12), S, Q(12));
       --Q14 : MUX4S port map (I1(13), I2(13), I3(13), I4(13), I5(13), I6(13), I7(13), I8(13), I9(13), I10(13), I11(13), I12(13), I13(13), I14(13), I15(13), I16(13), S, Q(13));
       --Q15 : MUX4S port map (I1(14), I2(14), I3(14), I4(14), I5(14), I6(14), I7(14), I8(14), I9(14), I10(14), I11(14), I12(14), I13(14), I14(14), I15(14), I16(14), S, Q(14));
       --Q16 : MUX4S port map (I1(15), I2(15), I3(15), I4(15), I5(15), I6(15), I7(15), I8(15), I9(15), I10(15), I11(15), I12(15), I13(15), I14(15), I15(15), I16(15), S, Q(15));
	

end ckt;