--==============================================================================================
--				LÓGICA DE UM MUX DE 2 BITS
--==============================================================================================
entity MUX2B is
	port (I : in bit_vector(1 downto 0);
			S : in bit_vector(1 downto 0);
			Y : out bit);
end MUX2B;

architecture ckt of MUX2B is

	begin

		Y <= (I(0) and (not S(1) and not S(0))) or (I(1) and (not S(1) and S(0)));

end ckt;

--==============================================================================================
--				LÓGICA DE UM DESLOCADOR <<1
--==============================================================================================

